----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Olivier Chaligne
-- 
-- Create Date: 02.02.2020 10:37:40
-- Design Name: 4 bit register using D fli flops
-- Module Name: Tutorial2_4 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity D_FF_4bit_reg is -- I/O Settings description
    Port ( clk : in STD_LOGIC; -- clock set as input
           d : in STD_LOGIC_VECTOR (3 DOWNTO 0); -- clock set as input
           ena : in STD_LOGIC; -- ena as an input
           rst : in STD_LOGIC; -- rst as an input
           q : out STD_LOGIC_VECTOR (3 DOWNTO 0)); -- q set as output
end D_FF_4bit_reg;

architecture Behavioral of D_FF_4bit_reg is -- description of D-Flip Flop
begin
    process(clk) -- run process for every rising edge of the clock.
    begin
        if rst = '1' then -- if reset triggered 
            q <= "0000"; --set outputs to 0
        elsif (clk' event and clk='1') Then -- if clock turns to high
            if ena = '1' then -- and enable is triggered
            q <= d; -- outputs q changed to d
            end if;
        end if;
    end process;
    
end Behavioral;


